`define DELAY 20
module alu32_testbench(); 
reg [31:0] A,B;
reg [2:0] S;
wire OF,Z;
wire [31:0] R;

alu32 alu_test(R,OF,Z,A,B,S);

initial begin
		//AND
A = 32'b01010111000000001010000000101110;
B = 32'b00101010100011100101000101100011;
S = 3'b000;
#`DELAY;
A = 32'b10101010101010101010101010101010;
B = 32'b01010101010101010101010101010101; 
S = 3'b000;
#`DELAY;
A = 32'b11110111000001101000010100100001;
B = 32'b10110001001000110101000101111010; 
S = 3'b000;
#`DELAY;
	//OR
A = 32'b01010111000000001010000000101110;
B = 32'b00101010100011100101000101100011;
S = 3'b001;
#`DELAY;
A = 32'b11010111001001001010000000001010;
B = 32'b10100110010001000010000101101001;
S = 3'b001;
#`DELAY;
A = 32'b11110111000001101000010100100001;
B = 32'b10110001001000110101000101111010; 
S = 3'b001;
#`DELAY;
		//ADDER
A = 32'b01000000000000000000000000000000;
B = 32'b01000000000000000000000000000000;
S = 3'b010;
#`DELAY;
A = 32'b11010111001001001010000000001010;
B = 32'b10100110010001000010000101101001; 
S = 3'b010;
#`DELAY;
A = 32'b11110111000001101000010100100001;
B = 32'b10110001001000110101000101111010; 
S = 3'b010;
#`DELAY;
		//XOR
A = 32'b01010111000000001010000000101110;
B = 32'b00101010100011100101000101100011;
S = 3'b011;
#`DELAY;
A = 32'b11010111001001001010000000001010;
B = 32'b10100110010001000010000101101001;
S = 3'b011;
#`DELAY;
A = 32'b11110111000001101000010100100001;
B = 32'b10110001001000110101000101111010; 
S = 3'b011;
#`DELAY;
		//SUBTRACTOR
A = 32'b11010111001001001010000000001010;
B = 32'b10100110010001000010000101101001;
S = 3'b100;
#`DELAY;
A = 32'b00000000000000000000000000100000;
B = 32'b00000000000000000000000000000010;
S = 3'b100;
#`DELAY;
A = 32'b00000000100100000000000001110000;
B = 32'b00000000000000001000000000000000;
#`DELAY;
		//ARITHMETIC RIGHT SHIFT
A = 32'b01010111000000001010000000101110;
B = 32'b00000000000000000000000000000001;
S = 3'b101;
#`DELAY;
A = 32'b11010111001001001010000000001010;
B = 32'b00000000000000000000000000000011; 
S = 3'b101;
#`DELAY;
A = 32'b11110111000001101000010100100001;
B = 32'b00000000000000000000000000001011;
S = 3'b101;
#`DELAY;
		//SHIFT LEFT
A = 32'b01010111000000001010000000101110;
B = 32'b00000000000000000000000000000001;
S = 3'b110;
#`DELAY;
A = 32'b11010111001001001010000000001010;
B = 32'b00000000000000000000000000000011; 
S = 3'b110;
#`DELAY;
A = 32'b11110111000001101000010100100001;
B = 32'b00000000000000000000000000001011;
S = 3'b110;
#`DELAY;
		//NOR
A = 32'b01010111000000001010000000101110;
B = 32'b00101010100011100101000101100011;
S = 3'b111;
#`DELAY;
A = 32'b11010111001001001010000000001010;
B = 32'b10100110010001000010000101101001;
S = 3'b111;
#`DELAY;
A = 32'b11110111000001101000010100100001;
B = 32'b10110001001000110101000101111010; 
S = 3'b111;
#`DELAY;
	
end
initial
begin
$monitor("time = %2d, Operation: %3b, A =%32b, B=%32b, R=%32b Owerflow=%1b, ZeroBit=%1b", $time, S,A, B, R,OF,Z);
end
 
endmodule